module controlador(input reset, input uart_redy,output en, output send_uart);
	
endmodule
